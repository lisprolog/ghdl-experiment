entity HalloWelt is
end entity;

architecture Verhalten of HalloWelt is
begin
	process
	begin
		-- Comment
		report "Hallo Welt";
		wait;
	end process;
end architecture;
