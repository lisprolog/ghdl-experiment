

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
PACKAGE MY IS
    FUNCTION INT_TO7SEG (A:INTEGER) RETURN STD_LOGIC_VECTOR;
	 PROCEDURE SEG_CTRL (SIGNAL NUMBER:IN INTEGER; SIGNAL DIGIT1,DIGIT2,DIGIT3,DIGIT4: OUT INTEGER RANGE 0 TO 9);
END MY;
 
 
PACKAGE BODY MY IS
   FUNCTION INT_TO7SEG (A:INTEGER) RETURN STD_LOGIC_VECTOR IS
	VARIABLE RESULT: STD_LOGIC_VECTOR(6 downto 0);
	BEGIN
	CASE A IS
	  WHEN 0 => RESULT:="1000000";
	  WHEN 1 => RESULT:="1111001";
	  WHEN 2 => RESULT:="0100100";
	  WHEN 3 => RESULT:="0110000";
	  WHEN 4 => RESULT:="0011001";
	  WHEN 5 => RESULT:="0010010";
	  WHEN 6 => RESULT:="0000010";
	  WHEN 7 => RESULT:="1111000";
	  WHEN 8 => RESULT:="0000000";
	  WHEN 9 => RESULT:="0010000";
	  WHEN OTHERS => RESULT:=(OTHERS=>'0');
	END CASE;
 
	RETURN RESULT;
	END INT_TO7SEG;
   --------------------------------------------------
	PROCEDURE SEG_CTRL (SIGNAL NUMBER:IN INTEGER; SIGNAL DIGIT1,DIGIT2,DIGIT3,DIGIT4: OUT INTEGER RANGE 0 TO 9) IS
	VARIABLE TEMP: INTEGER RANGE 0 TO 9999;
	VARIABLE D1: INTEGER RANGE 0 TO 9;
	VARIABLE D2: INTEGER RANGE 0 TO 9;
	VARIABLE D3: INTEGER RANGE 0 TO 9;
	VARIABLE D4: INTEGER RANGE 0 TO 9;
	BEGIN
	TEMP:=NUMBER;
	IF(TEMP>999)THEN
	 D4:=TEMP/1000;
	 TEMP:=TEMP-D4*1000;
	 ELSE
	 D4:=0;
	END IF;
	IF(TEMP>99)THEN
	 D3:=TEMP/100;
	 TEMP:=TEMP-D3*100;
	 ELSE
	 D3:=0;
	END IF;
	IF(TEMP>9)THEN
	 D2:=TEMP/10;
	 TEMP:=TEMP-D2*10;
	 ELSE
	 D2:=0;
	END IF;
	D1:=TEMP;
	DIGIT1<=D1;
	DIGIT2<=D2;
	DIGIT3<=D3;
	DIGIT4<=D4;
   END SEG_CTRL;
END MY;


